module segment7(in, negsigs);
    input[31:0] in;
    output[7:0] negsigs;

    wire[31:0] sigs;
    assign negsigs = ~sigs[7:0];
    mux32_32 MUX(sigs, in[4:0], {24'b0, 8'b11111101}, {24'b0, 8'b01100001}, {24'b0, 8'b11011011}, {24'b0, 8'b11110011}, {24'b0, 8'b01100111}, {24'b0, 8'b10110111}, {24'b0, 8'b10111111}, {24'b0, 8'b11100001}, {24'b0, 8'b11111111}, {24'b0, 8'b11100111}, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0, 32'b0);
endmodule